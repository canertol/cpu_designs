module INST_MEM (A,RD);
input [31:0] A;
output [31:0] RD;

reg [31:0] INST[88:0];

initial begin
 INST[0]  = 32'b1110_000_0010_0_1111_0000_0000_0000_1111; //	    SUB R0, R15, R15 	; R0 = 0
  INST[4] = 32'b1110_010_1100_0_0000_0000_0000_0000_0000; //		 STR  R0, R0 	      ; R0 = 0
 INST[8] = 32'b1110_010_1100_1_0000_0001_0000_0000_0000; //		    LDR R1, [R0, #0] 	; R1 = 0
  
 INST[12]  = 32'b1110_001_0100_0_0000_0010_0000_0000_0101; // 		 ADD R2, R0, #5 		; R2 = 5
 
 INST[16]  = 32'b1110_001_0100_0_0010_0011_0000_0000_0111; // 		 ADD R3, R2, #7		; R3 = R2 + 7 = 12
   INST[20] = 32'b1110_010_1100_0_0000_0011_0000_0000_0001; //		 STR  R3, [R0, #1] 	; R0 = 0
 INST[24] = 32'b1110_010_1100_1_0000_0001_0000_0000_0001; //		 LDR R1, [R0, #1] 	; R1 = 12  // 7ND inst
 
 
 INST[28] = 32'b1110_001_0010_0_0011_0111_0000_0000_1001; // 		 SUB R7, R3, #9 		; R7 = 3
 
 INST[32] = 32'b1110_000_1100_0_0111_0100_0000_0000_0010; // 		 ORR R4, R7, R2 		; R4 = 3 OR 5 = 7
 INST[36] = 32'b1110_010_1100_0_0000_0100_0000_0000_0111; //		 STR R4, [R0, #7] 	; R4 = 7
 INST[40] = 32'b1110_010_1100_1_0000_0001_0000_0000_0111; //		 LDR R1, [R0, #7] 	; R1 = 7 // 11ND inst
 
 INST[44] = 32'b1110_000_0000_0_0011_0101_0000_0000_0100; // 		 AND R5, R3, R4 		; R5 = 12 AND 7 = 4
 INST[48] = 32'b1110_010_1100_0_0000_0101_0000_0000_0011; //		 STR R5, [R0, #3] 	; R5 = 4
 INST[52] = 32'b1110_010_1100_1_0000_0001_0000_0000_0011; //		 LDR R1, [R0, #3] 	; R1 = 4  // 14ND inst
 
 INST[56] = 32'b1110_000_1101_0_0000_0010_00001_01_0_0001; //		 LSR  R2, R1, #1
 INST[60] = 32'b1110_010_1100_0_0000_0010_0000_0000_0100; //		 STR R2, [R0, #4] 	; R2 = 2
 INST[64] = 32'b1110_010_1100_1_0000_0001_0000_0000_0100; //		 LDR R1, [R0, #4] 	; R1 = 2   // 17ND inst
 
 
 INST[68] = 32'b1110_000_1010_1_0001_0000_0000_0000_0010;//			 CMP R1, R2
 
 INST[72] = 32'b1110_000_0100_0_1111_1111_0000_0000_0000; //		 ADD R15, R15, R0 	; PC = PC+8 (skips next)
 INST[76] = 32'b1110_001_0100_0_0000_0010_0000_0000_0001; //		 ADD R2, R0, #10 		; shouldn't happen
 
 INST[80] = 32'b1110_000_1101_0_0000_0010_00011_00_0_0010; //		 LSL  R2, #3  			; R2 = 16
  INST[84] = 32'b1110_010_1100_0_0000_0010_0000_0000_0101; //		 STR R2, [R0, #5] 	; R2 = 16
 INST[88] = 32'b1110_010_1100_1_0000_0010_0000_0000_0101; //		 LDR R2, [R0, #5] 	; R2 = 16
end 

assign RD = INST[A];

endmodule