module mux4_tb();
	reg [1:0] select;
	reg[3:0] mux_in1, mux_in2, mux_in3, mux_in4;
	wire [3:0] mux_out;
	reg[17:0] testvectors[63:0]; // array of testvectors
	reg [5:0] vectornum;

	mux4 #4 DUT(select, mux_in1,mux_in2,mux_in3,mux_in4, mux_out );
	
	// load vectors
	initial
	begin
	$readmemb("C:/Users/Caner/Documents/GitHub/Course-Projects/EE446/LAB1/mux4_tb.tv",testvectors);
	vectornum = 0;
	end
	
	//apply test vectors
	always
	begin
	 #5;
	 {mux_in1,mux_in2,mux_in3,mux_in4, select} = testvectors[vectornum];
	 vectornum = vectornum +1;
	end

endmodule
